localparam IDLE = 8'b00000000;//00
localparam START = 8'b00000001;//01
localparam ADDRESS = 8'b00000010;//02
localparam READ_ACK = 8'b00000100;//04
localparam WRITE_DATA = 8'b00001000;//08
localparam READ_DATA = 8'b00010000;//10
localparam READ_ACK2 = 8'b00100000;//20
localparam WRITE_ACK2 = 8'b01000000;//40
localparam STOP = 8'b10000000;//80
