localparam IDLE = 8'b00000000;
localparam START = 8'b00000001;
localparam ADDRESS = 8'b00000010;
localparam READ_ACK = 8'b00000100;
localparam WRITE_DATA = 8'b00001000;
localparam READ_DATA = 8'b00010000;
localparam READ_ACK2 = 8'b00100000;
localparam WRITE_ACK2 = 8'b01000000;
localparam STOP = 8'b10000000;
